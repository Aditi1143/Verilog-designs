module full_adder(a,b,cin,sum,cout);
input a,b,cin;
output sum,cout;
assign sum=a^b^cin;
assign cout=(a&b)|(cin&(a^b));
endmodule

module rca(a,b,cin,s,cout);
  input [3:0]a,b;
input cin;
output [3:0] s;
output cout;
  wire c1,c2,c3;
  full_adder f1(a[0],b[0],cin,s[0],c1);
  full_adder f2(a[1],b[1],c1,s[1],c2);
  full_adder f3(a[2],b[2],c2,s[2],c3);
  full_adder f4(a[3],b[3],c3,s[3],cout);
endmodule